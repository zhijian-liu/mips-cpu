`include "cpu/cpu.v"

module sopc(
	input	wire		clock,
	input	wire		reset
);

endmodule