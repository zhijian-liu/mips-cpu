module stage_wb(

);

endmodule