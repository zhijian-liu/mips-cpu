module cpu(
);